module Processor(
    input logic clock, reset
);

//Jazoolee//


//Thisara//


//Yasiru//



endmodule